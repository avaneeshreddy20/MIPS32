library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity dmem is
  port(
    memWrite,clk  : in std_logic;
    memRead       : in std_logic;
    address       : in std_logic_vector(9 downto 0);
    writeData     : in std_logic_vector(31 downto 0);
    readData      : out std_logic_vector(31 downto 0)
  );
end dmem;

architecture behavioral of dmem is
  signal readData1      : std_logic_vector(31 downto 0);
  type vector_of_mem is array(0 to 31) of std_logic_vector (31 downto 0);
  signal memory : vector_of_mem := ( 
        "00000000000000000000010101000000", 
        "00000011100000001011111100000101", 
        "00000000000000000000110000000000", 
        "00000000000000000100000000000000", 
        "00000000000000000000000000000011", 
        "00000000000000000000000000000111", 
        "00000000000000000000000000001111",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000"
    );
  begin
  
  readData <= memory(to_integer(unsigned(address))) when memRead = '1' else X"00000000";
  operationToDo : process(memWrite, address, writeData)
    begin

          if memWrite = '1' then
            memory(to_integer(unsigned(address))) <= writeData;
          end if;
 
  end process operationToDo;
end behavioral;
